----------------------------------------------------------------
-- Copyright 2020 University of Alberta

-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at

--     http://www.apache.org/licenses/LICENSE-2.0

-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.vnir;

package img_buffer_pkg is
    --Generating 10 buffers for each, allowing for storage of up to 10 rows
    constant NUM_SWIR_ROW_FIFO : integer := 1;
    constant NUM_VNIR_ROW_FIFO : integer := 1;

    --Number of bits in swir and vnir fifo
    --chosen to be 80 because it can fill whole multiples of vnir and swir pixels (10 and 16 bits respectively)
    --this is the lpm_numwords parameter for scfifo. usually must be 2^x but I think this is fine when not using the 
    --usedw port
    constant FIFO_WORD_LENGTH : integer := 80;  

    --Number of words in swir and vnir fifo
    constant VNIR_FIFO_DEPTH : integer := 256;
    constant SWIR_FIFO_DEPTH : integer := 64;

    --imaging buffer vnir fifo words (pipeline stage 1)
    constant pixels_per_row   : integer := FIFO_WORD_LENGTH/vnir.PIXEL_BITS; --80/10 = 8

    subtype vnir_fifo_pixel is std_logic_vector(vnir.PIXEL_BITS-1 downto 0);
    type vnir_fifo_row is array (0 to pixels_per_row-1) of vnir_fifo_pixel;
    type vnir_fifo_array is array (0 to VNIR_FIFO_DEPTH-1) of vnir_fifo_row;

    --vnir & swir row fragments are split into their respective FIFO word lengths
    subtype row_fragment_t is std_logic_vector (FIFO_WORD_LENGTH-1 downto 0);

    --The links between the vnir and swir fifos
    type vnir_link_a is array (0 to NUM_VNIR_ROW_FIFO-1) of row_fragment_t;
    type swir_link_a is array (0 to NUM_SWIR_ROW_FIFO-1) of row_fragment_t;

    type vnir_row_fragment_a is array (0 to VNIR_FIFO_DEPTH-1) of row_fragment_t;
    type swir_row_fragment_a is array (0 to SWIR_FIFO_DEPTH-1) of row_fragment_t;

    type row_type_buffer_a is array (0 to NUM_VNIR_ROW_FIFO-1) of vnir.row_type_t;

    
end package img_buffer_pkg;
